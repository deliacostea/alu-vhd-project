----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/12/2023 05:27:44 PM
-- Design Name: 
-- Module Name: wallace - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity wallace is
  Port (x, y: in std_logic_vector(31 downto 0);
  produs: out std_logic_vector(127 downto 0)
  
   );
end wallace;

architecture Behavioral of wallace is

component csa is
 Port ( a : in STD_LOGIC_VECTOR (63 downto 0);
        b : in STD_LOGIC_VECTOR (63 downto 0);
        c : in STD_LOGIC_VECTOR (63 downto 0);
        sum : out STD_LOGIC_VECTOR (63 downto 0);
        carry : out STD_LOGIC_VECTOR (63 downto 0));
end component;
signal x1,x2,x3,x4,x5,x6,x7,x8,x9,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20: std_logic_vector(63 downto 0) := (others => '0');
signal x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31,x32,x33,x34,x35,x36,x37,x38,x39,x40: std_logic_vector(63 downto 0):= (others => '0');
signal x41,x42,x43,x44,x45,x46,x47,x48,x49,x50,x51,x52,x53,x54,x55,x56,x57,x58,x59,x60,x61,x62,x63,x64:std_logic_vector(63 downto 0):= (others => '0');
signal c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32:std_logic_vector(63 downto 0):= (others => '0');
signal c33,c34,c35,c36,c37,c38,c39,c40,c41,c42,c43,c44,c45,c46,c47,c48,c49,c50,c51,c52,c53,c54,c55,c56,c57,c58,c59,c60,c61,c62:std_logic_vector(63 downto 0):= (others => '0');
signal s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29,s30,s31,s32:std_logic_vector(63 downto 0):= (others => '0');
signal s33,s34,s35,s36,s37,s38,s39,s40,s41,s42,s43,s44,s45,s46,s47,s48,s49,s50,s51,s52,s53,s54,s55,s56,s57,s58,s59,s60,s61,s62:std_logic_vector(63 downto 0):= (others => '0');
signal aux:std_logic_vector(63 downto 0) := (others => '0');
signal b:std_logic_vector(63 downto 0):= (others => '0');
signal Com2: std_logic_vector(127 downto 0):= (others => '0');
signal produs2: std_logic_vector(127 downto 0):= (others => '0');
signal aux2,aux3: std_logic_vector(31 downto 0) := (others => '0');


begin

process(produs2)
begin
if (x(31) xor y(31)) = '1' then
produs<= (not produs2) + 1;
else produs<=produs2;
end if;
end process;

process(x,y)
begin
if x(31)='1' then
aux2<= (not x) +1;
else aux2<= x;
end if;
if y(31)='1' then
aux3<=(not y) +1;
else aux3<= y;
end if;
end process;


aux<=x"00000000"&aux2;
b<=x"00000000"&aux3;
x1 <= aux and(b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     &b(0)& b(0) &b(0)& b(0) &b(0)& b(0)& b(0)& b(0)
     );
x2 <= (aux(62 downto 0)&'0') and 
    (b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    &b(1)& b(1) &b(1)& b(1) &b(1)& b(1)& b(1)& b(1)
    );
x3 <= (aux(61 downto 0)&"00") and
      (b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) &
      b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) &
      b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) &
      b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2)
      & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) &
       b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) &
       b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2)
       &b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2) & b(2)

      );

x4 <= (aux(60 downto 0)&"000") and( b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) &
      b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) &
      b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) &
      b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3)
      &b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) &
       b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) &
        b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3)
        &b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) & b(3) 
            );

x5 <= (aux(59 downto 0)&"0000") and (b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) &
             b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4) & b(4));

x6 <= (aux(58 downto 0)&"00000") and(b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) &
              b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5) & b(5));

x7 <= (aux(57 downto 0)&"000000") and (b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) &
               b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6) & b(6));

x8 <= (aux(56 downto 0)&"0000000") and (b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) &
                b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7) & b(7));

x9 <= (aux(55 downto 0)&"00000000") and (b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) &
                 b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8) & b(8))
;

x10 <= (aux(54 downto 0)&"000000000") and (b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) &
 b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9) & b(9))
;

x11 <= (aux(53 downto 0)&"0000000000") and (b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) &
 b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10) & b(10))
;

x12 <= (aux(52 downto 0)&"00000000000") and (b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) &
 b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11) & b(11))
;

x13 <= (aux(51 downto 0)&"000000000000") and (b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
  b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) &
 b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12) & b(12))
;

x14 <= (aux(50 downto 0)&"0000000000000") and (b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) &
 b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13) & b(13))
;

x15 <= (aux(49 downto 0)&"00000000000000") and (b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
  b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) &
 b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14) & b(14))
;

x16 <= (aux(48 downto 0)&"000000000000000") and (b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
  b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) &
 b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15) & b(15))
;

x17 <= (aux(47 downto 0)&"0000000000000000") and (b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) &
 b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16) & b(16))
;

x18 <= (aux(46 downto 0)&"00000000000000000") and (b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
  b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) &
 b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17) & b(17))
;

x19 <= (aux(45 downto 0)&"000000000000000000") and (b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
  b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) &
 b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18) & b(18))
;

x20 <= (aux(44 downto 0)&"0000000000000000000") and (b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
  b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) &
 b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19) & b(19))
;

x21 <= (aux(43 downto 0)&"00000000000000000000") and (b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
  b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) &
 b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20) & b(20)
);

x22 <= (aux(42 downto 0)&"000000000000000000000") and (b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
  b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) &
 b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21) & b(21))
;

x23 <= (aux(41 downto 0)&"0000000000000000000000") and (b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) &
 b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22) & b(22))
;

x24 <= (aux(40 downto 0)&"00000000000000000000000") and (b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
  b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) &
 b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23) & b(23))
;
       
x25 <= (aux(39 downto 0)&"000000000000000000000000") and (b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
  b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) &
 b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24) & b(24))
;
       
x26 <= (aux(38 downto 0)&"0000000000000000000000000") and (b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
  b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) &
 b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25) & b(25))
;
       
x27 <= (aux(37 downto 0)&"00000000000000000000000000") and (b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) &
 b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26) & b(26))
;
       
 x28 <= (aux(36 downto 0)&"000000000000000000000000000") and (b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
  b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) &
 b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27) & b(27))
;
       
x29 <= (aux(35 downto 0)&"0000000000000000000000000000") and (b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
  b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) &
 b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28) & b(28))
;
       
 x30 <= (aux(34 downto 0)&"00000000000000000000000000000") and (b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
  b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) &
 b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29) & b(29))
;
       
 x31 <= (aux(33 downto 0)&"000000000000000000000000000000") and (b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) &
 b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30) & b(30))
;
       
x32 <= (aux(32 downto 0)&"0000000000000000000000000000000") and (b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) &
 b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31) & b(31))
;

x33 <=(others => '0'); --inmultirea cu 0
x34 <=(others => '0');   
x35 <=(others => '0');  
x36 <=(others => '0');   
x37 <=(others => '0');          
x38 <=(others => '0');
x39 <=(others => '0');
x40 <=(others => '0');
x41 <=(others => '0');   
x42 <=(others => '0'); 
x43 <=(others => '0');
x44 <=(others => '0');
x45 <=(others => '0'); 
x46 <=(others => '0'); 
x47 <=(others => '0');  
x48 <=(others => '0');
x49 <=(others => '0');
x50 <=(others => '0');
x51 <=(others => '0'); 
x52 <=(others => '0');     
x53 <=(others => '0');
x54 <=(others => '0');    
x55 <=(others => '0');
x56 <=(others => '0');
x57 <=(others => '0');
x58 <=(others => '0');
x59 <=(others => '0');
x60 <=(others => '0');
x61 <=(others => '0');
x62 <=(others => '0');
x63 <=(others => '0'); 
x64 <= (others => '0');

--nivel 1

csa1: csa port map(x1,x2,x3,s1,c1);
csa2: csa port map(x4,x5,x6,s2,c2);
csa3: csa port map(x7,x8,x9,s3,c3);
csa4: csa port map(x10,x11,x12,s4,c4);
csa5: csa port map(x13,x14,x15,s5,c5);
csa6: csa port map(x16,x17,x18,s6,c6);
csa7: csa port map(x19,x20,x21,s7,c7);
csa8: csa port map(x22,x23,x24,s8,c8);
csa9: csa port map(x25,x26,x27,s9,c9);
csa10: csa port map(x28,x29,x30,s10,c10);
csa11: csa port map(x31,x32,x33,s11,c11);
csa12: csa port map(x34,x35,x36,s12,c12);
csa13: csa port map(x37,x38,x39,s13,c13);
csa14: csa port map(x40,x41,x42,s14,c14);
csa15: csa port map(x43,x44,x45,s15,c15);
csa16: csa port map(x46,x47,x48,s16,c16);
csa17: csa port map(x49,x50,x51,s17,c17);
csa18: csa port map(x52,x53,x54,s18,c18);
csa19: csa port map(x55,x56,x57,s19,c19);
csa20: csa port map(x58,x59,x60,s20,c20);
csa21: csa port map(x61,x62,x63,s21,c21);

--nivel 2

csa22: csa port map(s1,c1,s2,s22,c22);
csa23: csa port map(c2,s3,c3,s23,c23);
csa24: csa port map(s4,c4,s5,s24,c24);
csa25: csa port map(c5,s6,c6,s25,c25);
csa26: csa port map(s7,c7,s8,s26,c26);
csa27: csa port map(c8,s9,c9,s27,c27);
csa28: csa port map(s10,c10,s11,s28,c28);
csa29: csa port map(c11,s12,c12,s29,c29);
csa30: csa port map(s13,c13,s14,s30,c30);
csa31: csa port map(c14,s15,c15,s31,c31);
csa32: csa port map(s16,c16,s17,s32,c32);
csa33: csa port map(c17,s18,c18,s33,c33);
csa34: csa port map(s19,c19,s20,s34,c34);
csa35: csa port map(c20,s21,c21,s35,c35);

--nivel 3
csa36: csa port map(s22,c22,s23,s36,c36);
csa37: csa port map(c23,s24,c24,s37,c37);
csa38: csa port map(s25,c25,s26,s38,c38);
csa39: csa port map(c26,s27,c27,s39,c39);
csa40: csa port map(s28,c28,s29,s40,c40);
csa41: csa port map(c29,s30,c30,s41,c41);
csa42: csa port map(s31,c31,s32,s42,c42);
csa43: csa port map(c32,s33,c33,s43,c43);
csa44: csa port map(s34,c34,s35,s44,c44);

--nivel 4

csa45: csa port map(s36,c36,s37,s45,c45);
csa46: csa port map(c37,s38,c38,s46,c46);
csa47: csa port map(s39,c39,s40,s47,c47);
csa48: csa port map(c40,s41,c41,s48,c48);
csa49: csa port map(s42,c42,s43,s49,c49);
csa50: csa port map(c43,s44,c44,s50,c50);

--nivel 5

csa51: csa port map(s45,c45,s46,s51,c51);
csa52: csa port map(c46,s47,c47,s52,c52);
csa53: csa port map(s48,c48,s49,s53,c53);
css54: csa port map(c49,s50,c50,s54,c54);

--nivel 6

csa55: csa port map(s51,c51,s52,s55,c55);
csa56: csa port map(c52,s53,c53,s56,c56);
csa57: csa port map(s54,c54,c35,s57,c57);

--nivel 7

csa58: csa port map(s55,c55,s56,s58,c58);
csa59: csa port map(c56,s57,c57,s59,c59);

--nivel 8
csa60: csa port map(s58,c58,s59,s60,c60);

--nivel 9

csa61: csa port map(c59,s60,c60,s61,c61);

--nivel 10
csa62: csa port map(s61,c61,x"0000000000000000",s62,c62);









produs2(127 downto 64)<=c62;
produs2(63 downto 0)<=s62;


end Behavioral;
